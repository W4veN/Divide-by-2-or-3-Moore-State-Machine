-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition
-- Created on Tue Dec 29 17:27:18 2020

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Dividedby2or3 IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        y1 : OUT STD_LOGIC;
        y2 : OUT STD_LOGIC
    );
END Dividedby2or3;

ARCHITECTURE BEHAVIOR OF Dividedby2or3 IS
    TYPE type_fstate IS (A,B,C,D,E,F,G);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= A;
            y1 <= '0';
            y2 <= '0';
        ELSE
            y1 <= '0';
            y2 <= '0';
            CASE fstate IS
                WHEN A =>
                    IF ((x = '1')) THEN
                        reg_fstate <= B;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= A;
                    END IF;

                    IF (NOT((x = '1'))) THEN
                        y2 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        y2 <= '0';
                    END IF;

                    IF (NOT((x = '1'))) THEN
                        y1 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        y1 <= '0';
                    END IF;
                WHEN B =>
                    IF (NOT((x = '1'))) THEN
                        reg_fstate <= C;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= D;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= B;
                    END IF;
                WHEN C =>
                    IF (NOT((x = '1'))) THEN
                        reg_fstate <= E;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= C;
                    END IF;

                    IF (NOT((x = '1'))) THEN
                        y2 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        y2 <= '0';
                    END IF;
                WHEN D =>
                    IF (NOT((x = '1'))) THEN
                        reg_fstate <= F;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= G;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= D;
                    END IF;

                    IF ((x = '1')) THEN
                        y1 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        y1 <= '0';
                    END IF;
                WHEN E =>
                    IF ((x = '1')) THEN
                        reg_fstate <= B;
                    ELSIF (NOT((x = '1'))) THEN
                        reg_fstate <= A;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= E;
                    END IF;

                    IF (NOT((x = '1'))) THEN
                        y2 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        y2 <= '0';
                    END IF;
                WHEN F =>
                    IF ((x = '1')) THEN
                        reg_fstate <= B;
                    ELSIF (NOT((x = '1'))) THEN
                        reg_fstate <= E;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= F;
                    END IF;

                    IF (NOT((x = '1'))) THEN
                        y2 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        y2 <= '0';
                    END IF;

                    IF (NOT((x = '1'))) THEN
                        y1 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        y1 <= '0';
                    END IF;
                WHEN G =>
                    IF (NOT((x = '1'))) THEN
                        reg_fstate <= F;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= G;
                    END IF;
                WHEN OTHERS => 
                    y1 <= 'X';
                    y2 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
